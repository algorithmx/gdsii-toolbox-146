VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
UNITS DISTANCE MICRONS 1000 ;

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.14 ;
  WIDTH 0.06 ;
  THICKNESS 0.5 ;
END Metal1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.14 ;
  WIDTH 0.06 ;
  THICKNESS 0.5 ;
END Metal2

LAYER Via1
  TYPE CUT ;
  SPACING 0.08 ;
END Via1
